`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:52:07 04/07/2025 
// Design Name: 
// Module Name:    barrel_shifter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module barrel_shifter (input [15:0]a, input [3:0]s, input lr, output [15:0]x);
 wire x1l, x1r, x2l, x2r, x3l, x3r, x4l, x4r, x5l, x5r, x6l, x6r, x7l, x7r, x8l, x8r, x9l, x9r, x10l, x10r,
x11l, x11r, x12l, x12r, x13l, x13r, x14l, x14r, x15l, x15r, x16l, x16r;

 // For left shift
 mux16_1 m1(a[15],1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,s,x1l);
 mux16_1 m2(a[14],a[15],1,1,1,1,1,1,1,1,1,1,1,1,1,1,s,x2l);
 mux16_1 m3(a[13],a[14],a[15],1,1,1,1,1,1,1,1,1,1,1,1,1,s,x3l);
 mux16_1 m4(a[12],a[13],a[14],a[15],1,1,1,1,1,1,1,1,1,1,1,1,s,x4l);
 mux16_1 m5(a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,1,1,1,1,1,1,s,x5l);
 mux16_1 m6(a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,1,1,1,1,1,s,x6l);
 mux16_1 m7(a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,1,1,1,1,s,x7l);
 mux16_1 m8(a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,1,1,1,s,x8l);
 mux16_1 m9(a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,1,1,s,x9l);
 mux16_1 m10(a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,1,s,x10l);
 mux16_1 m11(a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,1,s,x11l);
 mux16_1 m12(a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,1,s,x12l);
 mux16_1 m13(a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,1,s,x13l);
 mux16_1 m14(a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,1,s,x14l);
 mux16_1 m15(a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],1,s,x15l);
 mux16_1
m16(a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],s,x16l);


 // For right shift
 mux16_1 m17(a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],s,x1r);
 mux16_1 m18(a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,s,x2r);
 mux16_1 m19(a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,s,x3r);
 mux16_1 m20(a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,s,x4r);
 mux16_1 m21(a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,s,x5r);
 mux16_1 m22(a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,s,x6r);
 mux16_1 m23(a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,1,s,x7r);
 mux16_1 m24(a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,1,1,s,x8r);
 mux16_1 m25(a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,1,1,1,s,x9r);
 mux16_1 m26(a[6],a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,1,1,1,1,s,x10r);
 mux16_1 m27(a[5],a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,1,1,1,1,1,s,x11r);
 mux16_1 m28(a[4],a[3],a[2],a[1],a[0],1,1,1,1,1,1,1,1,1,1,1,s,x12r);
 mux16_1 m29(a[3],a[2],a[1],a[0],1,1,1,1,1,1,1,1,1,1,1,1,s,x13r);
 mux16_1 m30(a[2],a[1],a[0],1,1,1,1,1,1,1,1,1,1,1,1,1,s,x14r);
 mux16_1 m31(a[1],a[0],1,1,1,1,1,1,1,1,1,1,1,1,1,1,s,x15r);
 mux16_1 m32(a[0],1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,s,x16r);
 mux_2_1 m33(x1l, x1r, lr, x[15]);
 mux_2_1 m34(x2l, x2r, lr, x[14]);
 mux_2_1 m35(x3l, x3r, lr, x[13]);
 mux_2_1 m36(x4l, x4r, lr, x[12]);
 mux_2_1 m37(x5l, x5r, lr, x[11]);
 mux_2_1 m38(x6l, x6r, lr, x[10]);
 mux_2_1 m39(x7l, x7r, lr, x[9]);
 mux_2_1 m40(x8l, x8r, lr, x[8]);
 mux_2_1 m41(x9l, x9r, lr, x[7]);
 mux_2_1 m42(x10l, x10r, lr, x[6]);
 mux_2_1 m43(x11l, x11r, lr, x[5]);
 mux_2_1 m44(x12l, x12r, lr, x[4]);
 mux_2_1 m45(x13l, x13r, lr, x[3]);
 mux_2_1 m46(x14l, x14r, lr, x[2]);
 mux_2_1 m47(x15l, x15r, lr, x[1]);
 mux_2_1 m48(x16l, x16r, lr, x[0]);
endmodule
